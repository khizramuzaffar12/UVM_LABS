class ahb_txn extends uvm_sequence_item;

  rand bit        write;
  rand bit [31:0] addr;
  rand bit [31:0] data;

  constraint addr_align { addr[1:0] == 2'b00; }

  // --------------------------------------------------
  // Factory + Field Registration
  // --------------------------------------------------
  `uvm_object_utils_begin(ahb_txn)
    `uvm_field_int(write, UVM_ALL_ON)
    `uvm_field_int(addr,  UVM_ALL_ON)
    `uvm_field_int(data,  UVM_ALL_ON)
  `uvm_object_utils_end

  // --------------------------------------------------
  // Constructor
  // --------------------------------------------------
  function new(string name = "ahb_txn");
    super.new(name);
  endfunction

endclass


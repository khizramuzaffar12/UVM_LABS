package ahb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ahb_txn.sv"
  `include "ahb_sequencer.sv"
  `include "ahb_driver.sv"
  `include "ahb_monitor.sv"
  `include "ahb_agent.sv"
  `include "ahb_scoreboard.sv"
  `include "ahb_env.sv"
  `include "ahb_sequence.sv"
  `include "ahb_test.sv"
endpackage


`timescale 1ns/1ns
import uvm_pkg::*;

module tb_top;

  initial begin
    run_test();
  end

endmodule

